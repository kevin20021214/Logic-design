module stateTrasition(
	output wire [6:0] display,
	output wire [3:0] digit,
	output trig,
	input echo,
	inout wire PS2_DATA,
	inout wire PS2_CLK,
	input wire rst,
	input wire clk
	);

    wire clk_1hz;
    clock_divider #(.n(26)) clk1h(.clk(clk), .clk_div(clk_1hz));

    wire [19:0] distance;

    parameter START = 0;
    parameter PLAY = 1;
    parameter LOSE = 2;
    parameter WIN = 3;
    reg [1:0]state, next_state;

    reg [9:0] sec, next_sec;
    wire [15:0] nums;

    // board
    wire [511:0] key_down;
    wire [8:0] last_change;
    wire been_ready;
    reg [3:0] key_num;
    parameter [8:0] KEY_CODES [0:21] = {
    	9'b0_0100_0101,	// 0 => 45
    	9'b0_0001_0110,	// 1 => 16
    	9'b0_0001_1110,	// 2 => 1E
    	9'b0_0010_0110,	// 3 => 26
    	9'b0_0010_0101,	// 4 => 25
    	9'b0_0010_1110,	// 5 => 2E
    	9'b0_0011_0110,	// 6 => 36
    	9'b0_0011_1101,	// 7 => 3D
    	9'b0_0011_1110,	// 8 => 3E
    	9'b0_0100_0110,	// 9 => 46
    
    	9'b0_0111_0000, // right_0 => 70
    	9'b0_0110_1001, // right_1 => 69
    	9'b0_0111_0010, // right_2 => 72
    	9'b0_0111_1010, // right_3 => 7A
    	9'b0_0110_1011, // right_4 => 6B
    	9'b0_0111_0011, // right_5 => 73
    	9'b0_0111_0100, // right_6 => 74
    	9'b0_0110_1100, // right_7 => 6C
    	9'b0_0111_0101, // right_8 => 75
    	9'b0_0111_1101,  // right_9 => 7D

    	9'b0_0101_1010,//enter=>5A
    	9'b0_0010_1001//space=>29
    };
    bin2bcd a(
        .bin(sec),
        .bcd(nums)
    );
    sonic_top B(
    	.clk(clk), 
       .rst(rst), 
       .Echo(echo), 
       .Trig(trig),
       .distance(distance)
    );

    KeyboardDecoder key_de (
    	.key_down(key_down),
    	.last_change(last_change),
    	.key_valid(been_ready),
    	.PS2_DATA(PS2_DATA),
    	.PS2_CLK(PS2_CLK),
    	.rst(rst),
    	.clk(clk)
    );
    My_SevenSegment sv(
    	.display(display),
    	.digit(digit),
    	.nums(nums),
    	.rst(rst),
    	.clk(clk)
    );
    //sec
    always @(posedge clk_1hz or posedge rst_1pulse) begin
    	if(rst_1pulse) sec<=0;
    	else if(state==play) sec<=next_sec;
        else sec<=0;
    end
    always @(*) begin
    	if(state==play) next_sec=sec+1;
    	else next_sec=0;
    end
    //state
    always @(posedge clk or posedge rst_1pulse) begin
    	if(rst_1pulse) state<=start;
    	else begin
    		case (state)
            start:begin 
                if(been_ready && key_down[last_change] == 1 && key_num == 10) state<=play;
                else state <= state; 
            end
            play:begin
                if(sec >= 300) state <= lose;
    			else if(distance < 50) state <= win;
                else state <= state;
            end
            lose:begin
                if(been_ready&&key_down[last_change]==1&&key_num==10) state<=start;
                else state<=state;
            end
    		win:begin
    			if(been_ready&&key_down[last_change]==1&&key_num==10) state<=start;
                else state<=state;
    		end
    		default: next_state<=state;
    		endcase
        end
    end
    //led
    always @(posedge clk or posedge rst_1pulse) begin
    	if(rst_1pulse) LED<=0;
    	else LED<=next_led;
    end
    always @(*) begin
    	case (state)
        start:next_led=16'b0000000000000000;
        play:next_led=16'b0000000000000001;
        lose:next_led=16'b1111111111111111;
    	win:next_led=16'b0000000011111111;
        default:next_led=LED;
    	endcase
    end

    //key_of_keyboard
    always @ (*) begin
    	case (last_change)
    		KEY_CODES[00]: key_num = 4'b0000;
    		KEY_CODES[01]: key_num = 4'b0001;
    		KEY_CODES[02]: key_num = 4'b0010;
    		KEY_CODES[03]: key_num = 4'b0011;
    		KEY_CODES[04]: key_num = 4'b0100;
    		KEY_CODES[05]: key_num = 4'b0101;
    		KEY_CODES[06]: key_num = 4'b0110;
    		KEY_CODES[07]: key_num = 4'b0111;
    		KEY_CODES[08]: key_num = 4'b1000;
    		KEY_CODES[09]: key_num = 4'b1001;
    		KEY_CODES[10]: key_num = 4'b0000;
    		KEY_CODES[11]: key_num = 4'b0001;
    		KEY_CODES[12]: key_num = 4'b0010;
    		KEY_CODES[13]: key_num = 4'b0011;
    		KEY_CODES[14]: key_num = 4'b0100;
    		KEY_CODES[15]: key_num = 4'b0101;
    		KEY_CODES[16]: key_num = 4'b0110;
    		KEY_CODES[17]: key_num = 4'b0111;
    		KEY_CODES[18]: key_num = 4'b1000;
    		KEY_CODES[19]: key_num = 4'b1001;

    		KEY_CODES[20]:key_num=4'b1010;
    		KEY_CODES[21]:key_num=4'b1011;

    		default : key_num = 4'b1111;
    	endcase
    end
endmodule



module my_clock_divider #(parameter n = 28'd2)
(
    input clock_in,
    output reg clock_out
);
reg [27:0] counter = 28'd0;
always @(posedge clock_in) begin
    counter <= counter + 1;
    if(counter >= (n-1)) begin
        counter <= 0;
    end
    clock_out <= (counter < n/2) ? 1'b1 : 1'b0;
end
endmodule 

module My_SevenSegment(
	output reg [6:0] display,
	output reg [3:0] digit,
	input wire [15:0] nums,
	input wire rst,
	input wire clk
    );
    
    reg [15:0] clk_divider;
    reg [3:0] display_num;
    
    always @ (posedge clk, posedge rst) begin
    	if (rst) begin
    		clk_divider <= 15'b0;
    	end else begin
    		clk_divider <= clk_divider + 15'b1;
    	end
    end
    
    always @ (posedge clk_divider[15], posedge rst) begin
    	if (rst) begin
    		display_num <= 4'b0000;
    		digit <= 4'b1111;
    	end else begin
    		case (digit)
    			4'b1110 : begin
    					display_num <= nums[7:4];
    					digit <= 4'b1101;
    				end
    			4'b1101 : begin
						display_num <= nums[11:8];
						digit <= 4'b1011;
					end
    			4'b1011 : begin
						display_num <= nums[15:12];
						digit <= 4'b0111;
					end
    			4'b0111 : begin
						display_num <= nums[3:0];
						digit <= 4'b1110;
					end
    			default : begin
						display_num <= nums[3:0];
						digit <= 4'b1110;
					end				
    		endcase
    	end
    end
    
    always @ (*) begin
    	case (display_num)
    		0 : display = 7'b1000000;	//0000
			1 : display = 7'b1111001;   //0001                                                
			2 : display = 7'b0100100;   //0010                                                
			3 : display = 7'b0110000;   //0011                                             
			4 : display = 7'b0011001;   //0100                                               
			5 : display = 7'b0010010;   //0101                                               
			6 : display = 7'b0000010;   //0110
			7 : display = 7'b1111000;   //0111
			8 : display = 7'b0000000;   //1000
			9 : display = 7'b0010000;	//1001
			
			10:display=7'b0111111;//-
			default : display = 7'b1111111;
    	endcase
    end
    
endmodule

module clock_divider #(
    parameter n = 27
)(
    input wire  clk,
    output wire clk_div  
);

    reg [n-1:0] num;
    wire [n-1:0] next_num;

    always @(posedge clk) begin
        num <= next_num;
    end

    assign next_num = num + 1;
    assign clk_div = num[n-1];
endmodule

module bin2bcd (
    input [9:0] bin,
    output reg [15:0] bcd
);
    integer i;
    always @(bin) begin
    bcd = 0;		 	
    for(i=0; i<=9; i=i+1) begin
        if(bcd[3:0]>4) begin
            bcd[3:0] = bcd[3:0] + 3;
        end
        if(bcd[7:4]>4) begin
            bcd[7:4] = bcd[7:4] + 3;
        end
        if(bcd[11:8]>4) begin
            bcd[11:8] = bcd[11:8] + 3;
        end
        if(bcd[15:12]>4) begin
            bcd[15:12] = bcd[15:12] + 3;
        end
        bcd = {bcd[14:0], bin[9-i]};
    end
end
endmodule

module div(clk, out_clk);
    input clk;
    output out_clk;
    reg out_clk;
    reg [6:0]cnt;
    
    always @(posedge clk) begin   
        if(cnt < 7'd50) begin
            cnt <= cnt + 1'b1;
            out_clk <= 1'b1;
        end 
        else if(cnt < 7'd100) begin
	        cnt <= cnt + 1'b1;
	        out_clk <= 1'b0;
        end
        else if(cnt == 7'd100) begin
            cnt <= 0;
            out_clk <= 1'b1;
        end
    end
endmodule